module adder(sum,carry,a,b)
