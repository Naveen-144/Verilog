module testbench ( );

// Inputs
reg [2:0] a;
reg [3:0] b;

// Outputs
wire [6:0] out;


// Instantiate the Design Under Test (DUT)
 product dut (
.a(a),
.b(b),
.res(out)
);

  // Clock and reset signals
  reg clk;
  reg rst;

  // Initial values
  initial begin
    clk = 0;
    rst = 1;
    #20;
    rst = 0;
  end

  // Clock generator
  always begin
    #10 clk = ~clk;
  end

  // Test sequence
  reg [3:0] i;
  always @(posedge clk, posedge rst) begin
    if (rst) begin
      i = 0;
    end else begin
      // Apply all possible val values (0-9)
      a <= $random%8;
	  b <= $random%16;
      #20;
      i = i + 1;
      if (i == 10) $finish;
    end
     $monitor("%d: a = %b, b = %b, res = %b", $time, a, b, out);
  end 
endmodule